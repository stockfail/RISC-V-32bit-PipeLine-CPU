`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:2**8-1];

    initial begin
       // $readmemh("code.mem", rom);
    // DATA Hazard Test
    rom[0] = 32'b0000000_00001_00010_000_00100_0110011; // add x4,x2,x1 -> 11+12=23
    rom[1] = 32'b0100000_00001_00100_000_00101_0110011; // sub x5,x4,x1 -> 23-11=12 // EX hazard
    rom[2] = 32'b0000000_00101_00100_000_00110_0110011; // add x6,x4,x5 -> 23+12=35 // EX + MEM hazard
    // Load Use Data Hazard Test
    rom[3] = 32'b0000000_00010_00000_010_01000_0100011; // sw x2,8(x0)
    rom[4] = 32'b000000001000_00000_010_00111_0000011; // lw x7,8(x0)
    rom[5] = 32'b0000000_00111_00001_000_01000_0110011; // add x8,x1,x7 -> 11+12=23 // Load Use Data hazard
    rom[6] = 32'b0000000_00010_00010_000_01001_0110011; // add x9,x2,x2 -> 24 // MEM hazard
    // Control Hazard Test
    // Branch Not Taken
    rom[7]  = 32'b0000000_00100_00101_000_01010_1100011; // beq x4, x5, +8   (23!=12 -> not taken)
    rom[8]  = 32'b0000000_00001_00010_000_01010_0110011; // add x10, x2, x1   (12+11=23, 실행됨)
    rom[9]  = 32'b0000000_00010_00001_000_01011_0110011; // add x11, x1, x2   (11+12=23, 실행됨)

    // Branch Taken (flush 1 instruction)
    rom[10] = 32'b0000000_00001_00001_000_01100_1100011; // beq x1, x1, +12  (taken, target=PC+12 → rom[13])
    rom[11] = 32'b0000000_00010_00001_000_01100_0110011; // add x12, x2, x1   (flush, 실행X) // hazard
    rom[12] = 32'b0000000_00010_00010_000_01101_0110011; // add x13, x2, x2   (jump, 실행X) // hazard
    rom[13] = 32'b0000000_00001_00010_000_01110_0110011; // add x14, x2, x1   (정상 실행됨)

    // JAL Test (flush 1 instruction)
    rom[14] = 32'b0_0000000100_0_00000000_00011_1101111; // jal x3, +8 (target=PC+8 → rom[16])
    rom[15] = 32'b0000000_00001_00001_000_01111_0110011; // add x15, x1, x1 (flush, 실행X) // hazard
    rom[16] = 32'b0000000_00010_00010_000_10000_0110011; // add x16, x2, x2 (정상 실행) // hazard 2번 반복 예상
    rom[17] = 32'b0000000_00010_00010_000_10001_0110011; // add x17, x2, x2 (정상 실행)
    rom[18] = 32'b0000000_00001_00010_000_10010_0110011; // add x18, x2, x1 (정상 실행)

    // JALR Test (flush 1 instruction)
    rom[19] = 32'b000001011000_00000_000_00011_1100111; // jalr x3, x0, +88 (target=88=rom[22])
    rom[20] = 32'b0000000_00001_00001_000_10011_0110011; // add x19, x1, x1 (flush, 실행X) // hazard
    rom[21] = 32'b0000000_00010_00010_000_10100_0110011; // add x20, x2, x2 (jump, 실행X) // hazard
    rom[22] = 32'b0000000_00001_00010_000_10101_0110011; // add x21, x2, x1 (정상 실행)
    end

    assign data = rom[addr[31:2]];
endmodule

/*
// Hazard Test
    rom[0] = 32'b0000000_00001_00010_000_00100_0110011; // add x4, x2, x1   (11+12=23)
    rom[1] = 32'b0100000_00001_00100_000_00101_0110011; // sub x5, x4, x1   (23-11=12)

    // Branch Not Taken
    rom[2] = 32'b0000000_00100_00101_000_00011_1100011; // beq x4, x5, +6   (23!=12 -> not taken)
    rom[3] = 32'b0000000_00001_00010_000_00110_0110011; // add x6, x2, x1   (12+11=23, 실행됨)
    rom[4] = 32'b0000000_00010_00001_000_00111_0110011; // add x7, x1, x2   (11+12=23, 실행됨)

    // Branch Taken (flush 1 instruction)
    rom[5] = 32'b0000000_00001_00001_000_01100_1100011; // beq x1, x1, +12  (target = 8) (11 == 11 -> taken -> 1 instruction flush)
    rom[6] = 32'b0000000_00001_00001_000_01000_0110011; // add x8, x1, x1   (flush, 실행X)
    rom[7] = 32'b0000000_00010_00010_000_01001_0110011; // add x9, x2, x2   (jump, 실행X) // Hazard 발생했다면 실행이됨
    rom[8] = 32'b0000000_00001_00010_000_01010_0110011; // add x10, x2, x1  (정상 실행됨)

    // JAL Test (flush 1 instruction)
   rom[9]  = 32'b0_0000000100_0_00000000_00011_1101111; // jal x3, +8 (target = 11)
   rom[10] = 32'b0000000_00001_00001_000_01011_0110011; // add x11, x1, x1 (flush, 실행X)
   rom[11] = 32'b0000000_00010_00010_000_01100_0110011; // add x12, x2, x2 (정상 실행)
   rom[12] = 32'b0000000_00010_00010_000_01101_0110011; // add x13, x2, x2 (정상 실행)
   rom[13] = 32'b0000000_00001_00010_000_01110_0110011; // add x14, x2, x1 (정상 실행)

    // JALR Test (flush 1 instruction)
    rom[14] = 32'b000001000100_00000_000_00011_1100111; // jalr x3, x0, +68 (target = 17)
    rom[15] = 32'b0000000_00001_00001_000_01111_0110011; // add x15, x1, x1 (flush, 실행X)
    rom[16] = 32'b0000000_00010_00010_000_10000_0110011; // add x16, x2, x2 (jump, 실행X)
    rom[17] = 32'b0000000_00001_00010_000_10001_0110011; // add x17, x2, x1 (정상 실행)
    //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // S-Type
    rom[18] = 32'b0000000_00010_00000_000_00011_0100011;// sb x2, 3(x0)
    rom[19] = 32'b0000000_00010_00000_001_00110_0100011;// sh x2, 6(x0)
    rom[20] = 32'b0000000_00010_00000_010_01000_0100011;// sw x2, 8(x0)
    //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // L-Type
    rom[21] = 32'b000000000011_00000_000_10010_0000011; // lb x18, 3(x0)
    rom[22] = 32'b000000000110_00000_001_10011_0000011; // lh x19, 6(x0)
    rom[23] = 32'b000000001000_00000_010_10100_0000011; // lw x20, 8(x0)
    rom[24] = 32'b000000000011_00000_100_10101_0000011; // lbu x21, 3(x0)
    rom[25] = 32'b000000000110_00000_101_10110_0000011; // lhu x22, 6(x0)
*/


 // rom[0] = 32'b0000000_00001_00010_000_00100_0110011;// add x4, x2, x1
    // rom[1] = 32'b0100000_00001_00100_000_00101_0110011;// sub x5, x4, x1
    // rom[2] = 32'b0000000_00010_00000_010_01000_0100011;// sw x2, 8(x0) 12를 메모리 저장
    // rom[3] = 32'b000000001000_00000_010_00110_0000011;// lw x6, 8(x0)  메모리에서 12값 x6에 로드
    // rom[4] = 32'b0000000_00001_00110_000_00111_0110011;// add x7, x6, x1
    // //rom[4] = 32'b0000000_00001_00010_000_00011_0110011;// add x3, x2, x1
    // rom[5] = 32'b0000000_00001_00110_000_01000_0110011;// add x8, x6, x1
    // rom[6] = 32'b
    //rom[x]=32'b fucn7 _ rs2 _ rs1 _f3 _ rd  _ op // R-Type
// rom[0] = 32'b0000000_00001_00010_000_00100_0110011;// add x4, x2, x1
// rom[1] = 32'b0100000_00001_00010_000_00101_0110011;// sub x5, x2, x1
// rom[2] = 32'b0000000_00000_00011_111_00110_0110011;// and x6, x3, x0
// rom[3] = 32'b0000000_00000_00011_110_00111_0110011;// or  x7, x3, x0
    //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // S-Type
//rom[4] = 32'b0000000_00010_00000_010_01000_0100011;// sw x2, 8(x0)
    //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // B-Type
//rom[5] = 32'b0000000_00010_00010_000_01100_1100011;// beq x2, x2, 12
    //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // L-Type
//rom[6] = 32'b000000001000_00000_010_01000_0000011;// lw x8, 8(x0)
    //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // I-Type
//rom[7] = 32'b000000000001_00001_000_01001_0010011;// addi x9, x1, 1 
//rom[8] = 32'b000000000100_00010_111_01010_0010011;// andi x10, x2, 4 
//rom[9] = 32'b000000000001_00010_110_01011_0010011;// ori x11, x2, 1 
//rom[10] = 32'b000000000011_00001_001_01100_0010011;// slli x12, x1, 1 // 2b00001011 << 3